/*
Program : 256x8-bit data memory (4-Byte blocks)
Author  : Isuru Nawinne
Date    : 30/05/2020

Description :

This program presents a primitive data memory module for CO224 Lab 6 - Part 2
This memory allows data to be read and written as 4-Byte blocks
*/
`timescale 1ns/100ps

module data_memory(
    clock,
    reset,
    read,
    write,
    address,
    writedata,
    readdata,
    busywait
);
input               clock;
input               reset;
input               read;
input               write;
input[5:0]          address;
input[31:0]         writedata;
output reg [31:0]   readdata;
output reg          busywait;

//Declare memory array 256x8-bits 
reg [7:0] memory_array [255:0];

//Detecting an incoming memory access
reg readaccess, writeaccess;
always @(read, write)
begin
    busywait = (read || write)? 1 : 0;
    readaccess = (read && !write)? 1 : 0;
    writeaccess = (!read && write)? 1 : 0;
end

//Reading & writing
always @(posedge clock)
begin
    if(readaccess)
    begin
        readdata[7:0]   = #40 memory_array[{address,2'b00}];
        readdata[15:8]  = #40 memory_array[{address,2'b01}];
        readdata[23:16] = #40 memory_array[{address,2'b10}];
        readdata[31:24] = #40 memory_array[{address,2'b11}];
        busywait = 0;
        readaccess = 0;
    end
    if(writeaccess)
    begin
        memory_array[{address,2'b00}] = #40 writedata[7:0];
        memory_array[{address,2'b01}] = #40 writedata[15:8];
        memory_array[{address,2'b10}] = #40 writedata[23:16];
        memory_array[{address,2'b11}] = #40 writedata[31:24];
        busywait = 0;
        writeaccess = 0;
    end
end

//Reset memory
integer i;
always @(posedge reset)
begin
    if (reset)
    begin
        for (i=0;i<256; i=i+1)
            memory_array[i] = 0;
        
        busywait = 0;
        readaccess = 0;
        writeaccess = 0;
    end
end

endmodule